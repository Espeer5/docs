--------------------------------------------------------------------------------
--                                                                            --
--  CORDIC16 Testbench                                                        --
--                                                                            --
--  This is atestbench for the CORDIC16 entity. It will test the CORDIC16     --
--  implementation architecture to ensure it can compute all desired          --
--  functions correctly over the appropriate range of input values. The       --
--  testbench entity is called CORDIC16_TB.                                   --
--                                                                            --
--  Revision History:                                                         --
--      12/5/2024  Edward Speer  Initial Revision                             --
--      12/6/2024  Edward Speer  Add test cases for all functions             --
--      12/8/2024  Edward Speer  Add full range of test vectors               --
--                                                                            --
--------------------------------------------------------------------------------

--
-- Imports
--

library ieee;
use     ieee.std_logic_1164.all;

entity CORDIC16_TB is
end    CORDIC16_TB;

--
-- CORDIC16_TB TB_architecture
--

architecture TB_architecture of CORDIC16_TB is

    --
    -- Component declaration of CORDIC16
    --

    component CORDIC16
        port (
            x : in  std_logic_vector(15 downto 0);  -- X input
            y : in  std_logic_vector(15 downto 0);  -- Y input
            f : in  std_logic_vector(4 downto 0);   -- Function selection signal
            r : out std_logic_vector(15 downto 0)   -- Result
        );
    end component;

    --
    -- Stimulus signals
    --

    signal x : std_logic_vector(15 downto 0);  -- X input
    signal y : std_logic_vector(15 downto 0);  -- Y input
    signal f : std_logic_vector(4 downto 0);   -- Function selection signal

    --
    -- Observed signals
    --

    signal r : std_logic_vector(15 downto 0);  -- Result

    --
    -- Test vectors
    --

    constant nTests : Integer := 44 * 4 + 2 * 40;
    signal   xs     : std_logic_vector(nTests * 16 - 1 downto 0);
    signal   ys     : std_logic_vector(nTests * 16 - 1 downto 0);
    signal   fs     : std_logic_vector(nTests * 5  - 1 downto 0);
    signal   rs     : std_logic_vector(nTests * 16 - 1 downto 0);

begin

    --
    -- Device under test port map
    --

    DUT : CORDIC16 port map (
        x => x,
        y => y,
        f => f,
        r => r
    );

    --
    -- Test vectors
    --
    ys <=   "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" & 
            "----------------" & 
            "----------------" & 
            "----------------" &
            "----------------" &
            "0000011001100110" &
            "0000100000000000" &
            "0000100110011010" &
            "0000101100110011" &
            "0000110011001101" &
            "0000111001100110" &
            "0001000000000000" &
            "0001000110011010" &
            "0001001100110011" &
            "0001010011001101" &
            "0001011001100110" &
            "0001100000000000" &
            "0001100110011010" &
            "0001101100110011" &
            "0001110011001101" &
            "0001111001100110" &
            "0010000000000000" &
            "0010000110011010" &
            "0010001100110011" &
            "0010010011001101" &
            "0010011001100110" &
            "0010100000000000" &
            "0010100110011010" &
            "0010101100110011" &
            "0010110011001101" &
            "0010111001100110" &
            "0011000000000000" &
            "0011000110011010" &
            "0011001100110011" &
            "0011010011001101" &
            "0011011001100110" &
            "0011100000000000" &
            "0011100110011010" &
            "0011101100110011" &
            "0011110011001101" &
            "0011111001100110" &
            "0100000000000000" &
            "0100000110011010" &
            "0100001100110011" &
            "0100010011001101" &
            "0000011001100110" &
            "0000100000000000" &
            "0000100110011010" &
            "0000101100110011" &
            "0000110011001101" &
            "0000111001100110" &
            "0001000000000000" &
            "0001000110011010" &
            "0001001100110011" &
            "0001010011001101" &
            "0001011001100110" &
            "0001100000000000" &
            "0001100110011010" &
            "0001101100110011" &
            "0001110011001101" &
            "0001111001100110" &
            "0010000000000000" &
            "0010000110011010" &
            "0010001100110011" &
            "0010010011001101" &
            "0010011001100110" &
            "0010100000000000" &
            "0010100110011010" &
            "0010101100110011" &
            "0010110011001101" &
            "0010111001100110" &
            "0011000000000000" &
            "0011000110011010" &
            "0011001100110011" &
            "0011010011001101" &
            "0011011001100110" &
            "0011100000000000" &
            "0011100110011010" &
            "0011101100110011" &
            "0011110011001101" &
            "0011111001100110" &
            "0100000000000000" &
            "0100000110011010" &
            "0100001100110011" &
            "0100010011001101";


    xs <=   "0000001000111100" &
            "0000010001111000" &
            "0000011010110100" &
            "0000100011110000" &
            "0000101100101100" &
            "0000110101100111" &
            "0000111110100011" &
            "0001000111011111" &
            "0001010000011011" &
            "0001011001010111" &
            "0001100010010011" &
            "0001101011001111" &
            "0001110100001011" &
            "0001111101000111" &
            "0010000110000011" &
            "0010001110111111" &
            "0010010111111010" &
            "0010100000110110" &
            "0010101001110010" &
            "0010110010101110" &
            "0010111011101010" &
            "0011000100100110" &
            "0011001101100010" &
            "0011010110011110" &
            "0011011111011010" &
            "0011101000010110" &
            "0011110001010010" &
            "0011111010001101" &
            "0100000011001001" &
            "0100001100000101" &
            "0100010101000001" &
            "0100011101111101" &
            "0100100110111001" &
            "0100101111110101" &
            "0100111000110001" &
            "0101000001101101" &
            "0101001010101001" &
            "0101010011100101" &
            "0101011100100000" &
            "0101100101011100" &
            "0101101110011000" &
            "0101110111010100" &
            "0110000000010000" &
            "0110001001001100" &
            "0000001000111100" &
            "0000010001111000" &
            "0000011010110100" &
            "0000100011110000" &
            "0000101100101100" &
            "0000110101100111" &
            "0000111110100011" &
            "0001000111011111" &
            "0001010000011011" &
            "0001011001010111" &
            "0001100010010011" &
            "0001101011001111" &
            "0001110100001011" &
            "0001111101000111" &
            "0010000110000011" &
            "0010001110111111" &
            "0010010111111010" &
            "0010100000110110" &
            "0010101001110010" &
            "0010110010101110" &
            "0010111011101010" &
            "0011000100100110" &
            "0011001101100010" &
            "0011010110011110" &
            "0011011111011010" &
            "0011101000010110" &
            "0011110001010010" &
            "0011111010001101" &
            "0100000011001001" &
            "0100001100000101" &
            "0100010101000001" &
            "0100011101111101" &
            "0100100110111001" &
            "0100101111110101" &
            "0100111000110001" &
            "0101000001101101" &
            "0101001010101001" &
            "0101010011100101" &
            "0101011100100000" &
            "0101100101011100" &
            "0101101110011000" &
            "0101110111010100" &
            "0110000000010000" &
            "0110001001001100" &
            "0000001000111100" &
            "0000010001111000" &
            "0000011010110100" &
            "0000100011110000" &
            "0000101100101100" &
            "0000110101100111" &
            "0000111110100011" &
            "0001000111011111" &
            "0001010000011011" &
            "0001011001010111" &
            "0001100010010011" &
            "0001101011001111" &
            "0001110100001011" &
            "0001111101000111" &
            "0010000110000011" &
            "0010001110111111" &
            "0010010111111010" &
            "0010100000110110" &
            "0010101001110010" &
            "0010110010101110" &
            "0010111011101010" &
            "0011000100100110" &
            "0011001101100010" &
            "0011010110011110" &
            "0011011111011010" &
            "0011101000010110" &
            "0011110001010010" &
            "0011111010001101" &
            "0100000011001001" &
            "0100001100000101" &
            "0100010101000001" &
            "0100011101111101" &
            "0100100110111001" &
            "0100101111110101" &
            "0100111000110001" &
            "0101000001101101" &
            "0101001010101001" &
            "0101010011100101" &
            "0101011100100000" &
            "0101100101011100" &
            "0101101110011000" &
            "0101110111010100" &
            "0110000000010000" &
            "0110001001001100" &
            "0000001000111100" &
            "0000010001111000" &
            "0000011010110100" &
            "0000100011110000" &
            "0000101100101100" &
            "0000110101100111" &
            "0000111110100011" &
            "0001000111011111" &
            "0001010000011011" &
            "0001011001010111" &
            "0001100010010011" &
            "0001101011001111" &
            "0001110100001011" &
            "0001111101000111" &
            "0010000110000011" &
            "0010001110111111" &
            "0010010111111010" &
            "0010100000110110" &
            "0010101001110010" &
            "0010110010101110" &
            "0010111011101010" &
            "0011000100100110" &
            "0011001101100010" &
            "0011010110011110" &
            "0011011111011010" &
            "0011101000010110" &
            "0011110001010010" &
            "0011111010001101" &
            "0100000011001001" &
            "0100001100000101" &
            "0100010101000001" &
            "0100011101111101" &
            "0100100110111001" &
            "0100101111110101" &
            "0100111000110001" &
            "0101000001101101" &
            "0101001010101001" &
            "0101010011100101" &
            "0101011100100000" &
            "0101100101011100" &
            "0101101110011000" &
            "0101110111010100" &
            "0110000000010000" &
            "0110001001001100" &
            "0100011001100110" &
            "0100010011001101" &
            "0100001100110011" &
            "0100000110011010" &
            "0100000000000000" &
            "0011111001100110" &
            "0011110011001101" &
            "0011101100110011" &
            "0011100110011010" &
            "0011100000000000" &
            "0011011001100110" &
            "0011010011001101" &
            "0011001100110011" &
            "0011000110011010" &
            "0011000000000000" &
            "0010111001100110" &
            "0010110011001101" &
            "0010101100110011" &
            "0010100110011010" &
            "0010100000000000" &
            "0010011001100110" &
            "0010010011001101" &
            "0010001100110011" &
            "0010000110011010" &
            "0010000000000000" &
            "0001111001100110" &
            "0001110011001101" &
            "0001101100110011" &
            "0001100110011010" &
            "0001100000000000" &
            "0001011001100110" &
            "0001010011001101" &
            "0001001100110011" &
            "0001000110011010" &
            "0001000000000000" &
            "0000111001100110" &
            "0000110011001101" &
            "0000101100110011" &
            "0000100110011010" &
            "0000100000000000" &
            "0100011001100110" &
            "0100010011001101" &
            "0100001100110011" &
            "0100000110011010" &
            "0100000000000000" &
            "0011111001100110" &
            "0011110011001101" &
            "0011101100110011" &
            "0011100110011010" &
            "0011100000000000" &
            "0011011001100110" &
            "0011010011001101" &
            "0011001100110011" &
            "0011000110011010" &
            "0011000000000000" &
            "0010111001100110" &
            "0010110011001101" &
            "0010101100110011" &
            "0010100110011010" &
            "0010100000000000" &
            "0010011001100110" &
            "0010010011001101" &
            "0010001100110011" &
            "0010000110011010" &
            "0010000000000000" &
            "0001111001100110" &
            "0001110011001101" &
            "0001101100110011" &
            "0001100110011010" &
            "0001100000000000" &
            "0001011001100110" &
            "0001010011001101" &
            "0001001100110011" &
            "0001000110011010" &
            "0001000000000000" &
            "0000111001100110" &
            "0000110011001101" &
            "0000101100110011" &
            "0000100110011010" &
            "0000100000000000";



    fs <=   "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00001" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00101" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00010" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00110" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "00100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100" &
            "01100";

    process      -- TEST_PROCESS
    begin

        -- Initialize DUT inputs
        x <= (others => '0');
        y <= (others => '0');
        f <= (others => '0');

        wait for 10 ns;

        -- Loop over test vectors and test each case
        for i in 0 to nTests - 1 loop
            x <= xs(i * 16 + 15 downto i * 16);
            y <= ys(i * 16 + 15 downto i * 16);
            f <= fs(i * 5  + 4  downto i * 5);

            wait for 10 ns;

            report std_logic'image(r(15)) & std_logic'image(r(14)) &
                   std_logic'image(r(13)) & std_logic'image(r(12)) &
                   std_logic'image(r(11)) & std_logic'image(r(10)) &
                   std_logic'image(r(9))  & std_logic'image(r(8))  &
                   std_logic'image(r(7))  & std_logic'image(r(6))  &
                   std_logic'image(r(5))  & std_logic'image(r(4))  &
                   std_logic'image(r(3))  & std_logic'image(r(2))  &
                   std_logic'image(r(1))  & std_logic'image(r(0))
                   severity note;
        end loop;

        -- End the simulation
        wait;

    end process; -- TEST_PROCESS


end TB_architecture;

configuration TESTBENCH_FOR_CORDIC16_IMPLEMENTATION of CORDIC16_TB is
    for TB_architecture
        for DUT : CORDIC16
            use entity work.CORDIC16(implementation);
        end for;
    end for;
end TESTBENCH_FOR_CORDIC16_IMPLEMENTATION;
