process (clk)
begin
    x <= a;
end process;